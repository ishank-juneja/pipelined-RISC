library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library std;
use std.standard.all;

entity decoder is
	port (t3 : in std_logic_vector(7 downto 0);
			input : in std_logic_vector(2 downto 0);
			next_t3 : out std_logic_vector(7 downto 0));
end entity;
architecture struct of decoder is
begin
	next_t3(0) <= t3(0) and not(not(input(2)) and not(input(1)) and not(input(0)));
	next_t3(1) <= t3(1) and not(not(input(2)) and not(input(1)) and     input(0))	;
	next_t3(2) <= t3(2) and not(not(input(2)) and     input(1)  and not(input(0)));
	next_t3(3) <= t3(3) and not(not(input(2)) and 	  input(1)  and 	  input(0))	;
	next_t3(4) <= t3(4) and not(	  input(2)  and not(input(1)) and not(input(0)));
	next_t3(5) <= t3(5) and not(	  input(2)  and not(input(1)) and 	  input(0))	;
	next_t3(6) <= t3(6) and not(	  input(2)  and 	  input(1)  and not(input(0)));
	next_t3(7) <= t3(7) and not(	  input(2)  and     input(1)  and 	  input(0))	;
end struct;